x"00d0",	--ladda in d0 till reg0
x"10d1",	--spara värdet i reg0 på d1
x"00d3",	--ladda in d3 till reg0
x"10d4", 	--spara värdet i reg0 på d4
x"00d1",	--ladda in värdet i d1 till reg0
x"20d3",	--addera reg0=reg0+d3
x"10d2",	--spara v'rdet i reg0 på d2	
x"02d1",	--ladda in det d1 pekar på till reg0
x"a2d2",	--jämför det värde d2 pekar på och värdet i reg0
x"b014",	--hoppa till adress 14 om resultat   det värdet d2 pekar på är större än det i reg0
x"00d2",	--ladda in d2 i reg0
x"10d1",	--spara värdet i reg0 på d1
x"a0d6",	--jämför det på reg0 och det i d6
x"c00f",	--beq, hoppa till f om det värde d6 pekar var större on det i reg0
x"6004",	--hoppa till adress 4
x"00d3",	--ladda in d3 på reg0
x"a0d4",	--cmp $d4 och reg0
x"c013",	--beq hoppa till 13 om $d4 var större än reg0
x"6000",	--hoppa till 00
x"8000",	--halt
x"02d1",	--ladda in det d1 pekar på till reg0
x"06d2",	--ladda in det d2 pekar till reg1
x"12d2",	--spara reg0 på den adress som d2 pekar
x"16d1",	--spara reg2 på den adress som d1 pekar på
x"00d5",	--ladda in d5 på reg0
x"10d4",	--spara värdet i reg0 på d4
x"600a",	--hoppa tll 10
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"00e0",
x"0000",
x"0000",
x"0001",
x"0000",
x"0000",
x"00ff",
x"0002",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"0000",
x"92f1",
x"8034",
x"971b",
x"99fb",
x"7ef1",
x"90e8",
x"5ee7",
x"3de3",
x"7351",
x"53ed",
x"56a2",
x"dea5",
x"6c5a",
x"835f",
x"7c67",
x"ec86",
x"bd89",
x"969c",
x"5f63",
x"72d7",
x"959f",
x"6081",
x"4c67",
x"7e12",
x"9fc4",
x"b11c",
x"623d",
x"8832",
x"78ea",
x"9f74",
x"7044",
x"bfb0",

