library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity pm is
	port (clk		: in std_logic;
		rst			: in std_logic;
		adress_pm	: in std_logic_vector(7 downto 0);
		pm_read		: in std_logic;
		pm_write	: in std_logic;
		bus_in		: in std_logic_vector(15 downto 0);
		bus_out		: out std_logic_vector(15 downto 0)
	);
end pm;

architecture Behavioral of pm is

	-- Declaration of a block-RAM with 256 addresses of 8 bits.
	type ram_t is array (0 to 255) of
	  std_logic_vector(15 downto 0);
	
	-- Original ram, used when reset button is used.
	signal original_ram : ram_t := (
		x"00ff",
		x"0812",
		x"f905",
		x"1812",
		x"600c",
		x"10f8",
		x"f90a",
		x"1812",
		x"00fe",
		x"600c",
		x"10f9",
		x"60a9",
		x"e000",
		x"0016",
		x"f111",
		x"1016",
		x"6013",
		x"d000",
		x"6000",
		x"00ff",
		x"20fe",
		x"a0fd",
		x"c000",
		x"6014",
		x"5106",
		x"14e0",
		x"20e0",
		x"5101",
		x"18e0",
		x"20e0",
		x"9000",
		x"1ce0",
		x"0cff",
		x"ace0",
		x"c000",
		x"20f6",
		x"9000",
		x"2cfe",
		x"6021",
		x"0022",
		x"f12f",
		x"1022",
		x"00f5",
		x"04f4",
		x"08ff",
		x"0cfb",
		x"6018",
		x"00f8",
		x"10f5",
		x"0422",
		x"f538",
		x"1422",
		x"04f4",
		x"08fe",
		x"0cfb",
		x"6018",
		x"0422",
		x"f540",
		x"1422",
		x"00f3",
		x"04f2",
		x"08ff",
		x"0cfb",
		x"6018",
		x"00f9",
		x"10f3",
		x"0422",
		x"f549",
		x"1422",
		x"04f2",
		x"08fe",
		x"0cfb",
		x"6018",
		x"00ed",
		x"5106",
		x"20ee",
		x"5101",
		x"9000",
		x"00e8",
		x"10ee",
		x"00e7",
		x"10ed",
		x"5106",
		x"20ee",
		x"5101",
		x"20fe",
		x"9000",
		x"00e2",
		x"9000",
		x"04e1",
		x"9400",
		x"0cfc",
		x"acff",
		x"c064",
		x"20fe",
		x"9000",
		x"acfe",
		x"c064",
		x"24fe",
		x"9400",
		x"00df",
		x"9000",
		x"04de",
		x"9400",
		x"0cfa",
		x"acff",
		x"c000",
		x"20fe",
		x"9000",
		x"acfe",
		x"c000",
		x"24fe",
		x"9400",
		x"6000",
		x"00ed",
		x"a0ff",
		x"c0a3",
		x"a0e4",
		x"c0a6",
		x"00ee",
		x"a0f7",
		x"c08d",
		x"a0f1",
		x"c07d",
		x"6027",
		x"00f3",
		x"a0ed",
		x"c0a0",
		x"20fe",
		x"a0ed",
		x"c0a0",
		x"20fe",
		x"a0ed",
		x"c0a0",
		x"20fe",
		x"a0ed",
		x"c0a0",
		x"00fc",
		x"20fe",
		x"10fc",
		x"60cc",
		x"00f5",
		x"a0ed",
		x"c09d",
		x"20fe",
		x"a0ed",
		x"c09d",
		x"20fe",
		x"a0ed",
		x"c09d",
		x"20fe",
		x"a0ed",
		x"c09d",
		x"00fa",
		x"20fe",
		x"10fa",
		x"60cc",
		x"00fe",
		x"10ec",
		x"607c",
		x"00ff",
		x"10ec",
		x"607c",
		x"00fe",
		x"10ea",
		x"6077",
		x"00ff",
		x"10ea",
		x"6077",
		x"00e6",
		x"a0eb",
		x"c0c1",
		x"00e5",
		x"a0e9",
		x"c0b6",
		x"00e6",
		x"20fe",
		x"10e6",
		x"00e5",
		x"20fe",
		x"10e5",
		x"6072",
		x"00ff",
		x"10e5",
		x"00ea",
		x"a0ff",
		x"00ed",
		x"c0be",
		x"20fe",
		x"60bf",
		x"30fe",
		x"10e7",
		x"60af",
		x"00ff",
		x"10e6",
		x"00ec",
		x"a0ff",
		x"00ee",
		x"c0c9",
		x"20fe",
		x"60ca",
		x"30fe",
		x"10e8",
		x"60ac",
		x"00f0",
		x"10e8",
		x"00ef",
		x"10e7",
		x"00f9",
		x"40fe",
		x"10ec",
		x"00fa",
		x"a0fb",
		x"c0da",
		x"00fc",
		x"a0fb",
		x"c0da",
		x"6027",
		x"00ff",
		x"10fa",
		x"10fc",
		x"6027",
		x"0050",
		x"0048",
		x"0000",
		x"0030",
		x"0038",
		x"0004",
		x"002e",
		x"0000",
		x"0000",
		x"0017",
		x"0020",
		x"0040",
		x"0000",
		x"0040",
		x"0000",
		x"0018",
		x"0020",
		x"0018",
		x"0020",
		x"003e",
		x"003f",
		x"0001",
		x"0002",
		x"0001",
		x"0080",
		x"0003",
		x"0000",
		x"0000",
		x"0000",
		x"0003",
		x"0000",
		x"0800",
		x"0001",
		x"0000"
	);
	
	--PM
	signal ram : ram_t := (
		x"00ff",
		x"0812",
		x"f905",
		x"1812",
		x"600c",
		x"10f8",
		x"f90a",
		x"1812",
		x"00fe",
		x"600c",
		x"10f9",
		x"60a9",
		x"e000",
		x"0016",
		x"f111",
		x"1016",
		x"6013",
		x"d000",
		x"6000",
		x"00ff",
		x"20fe",
		x"a0fd",
		x"c000",
		x"6014",
		x"5106",
		x"14e0",
		x"20e0",
		x"5101",
		x"18e0",
		x"20e0",
		x"9000",
		x"1ce0",
		x"0cff",
		x"ace0",
		x"c000",
		x"20f6",
		x"9000",
		x"2cfe",
		x"6021",
		x"0022",
		x"f12f",
		x"1022",
		x"00f5",
		x"04f4",
		x"08ff",
		x"0cfb",
		x"6018",
		x"00f8",
		x"10f5",
		x"0422",
		x"f538",
		x"1422",
		x"04f4",
		x"08fe",
		x"0cfb",
		x"6018",
		x"0422",
		x"f540",
		x"1422",
		x"00f3",
		x"04f2",
		x"08ff",
		x"0cfb",
		x"6018",
		x"00f9",
		x"10f3",
		x"0422",
		x"f549",
		x"1422",
		x"04f2",
		x"08fe",
		x"0cfb",
		x"6018",
		x"00ed",
		x"5106",
		x"20ee",
		x"5101",
		x"9000",
		x"00e8",
		x"10ee",
		x"00e7",
		x"10ed",
		x"5106",
		x"20ee",
		x"5101",
		x"20fe",
		x"9000",
		x"00e2",
		x"9000",
		x"04e1",
		x"9400",
		x"0cfc",
		x"acff",
		x"c064",
		x"20fe",
		x"9000",
		x"acfe",
		x"c064",
		x"24fe",
		x"9400",
		x"00df",
		x"9000",
		x"04de",
		x"9400",
		x"0cfa",
		x"acff",
		x"c000",
		x"20fe",
		x"9000",
		x"acfe",
		x"c000",
		x"24fe",
		x"9400",
		x"6000",
		x"00ed",
		x"a0ff",
		x"c0a3",
		x"a0e4",
		x"c0a6",
		x"00ee",
		x"a0f7",
		x"c08d",
		x"a0f1",
		x"c07d",
		x"6027",
		x"00f3",
		x"a0ed",
		x"c0a0",
		x"20fe",
		x"a0ed",
		x"c0a0",
		x"20fe",
		x"a0ed",
		x"c0a0",
		x"20fe",
		x"a0ed",
		x"c0a0",
		x"00fc",
		x"20fe",
		x"10fc",
		x"60cc",
		x"00f5",
		x"a0ed",
		x"c09d",
		x"20fe",
		x"a0ed",
		x"c09d",
		x"20fe",
		x"a0ed",
		x"c09d",
		x"20fe",
		x"a0ed",
		x"c09d",
		x"00fa",
		x"20fe",
		x"10fa",
		x"60cc",
		x"00fe",
		x"10ec",
		x"607c",
		x"00ff",
		x"10ec",
		x"607c",
		x"00fe",
		x"10ea",
		x"6077",
		x"00ff",
		x"10ea",
		x"6077",
		x"00e6",
		x"a0eb",
		x"c0c1",
		x"00e5",
		x"a0e9",
		x"c0b6",
		x"00e6",
		x"20fe",
		x"10e6",
		x"00e5",
		x"20fe",
		x"10e5",
		x"6072",
		x"00ff",
		x"10e5",
		x"00ea",
		x"a0ff",
		x"00ed",
		x"c0be",
		x"20fe",
		x"60bf",
		x"30fe",
		x"10e7",
		x"60af",
		x"00ff",
		x"10e6",
		x"00ec",
		x"a0ff",
		x"00ee",
		x"c0c9",
		x"20fe",
		x"60ca",
		x"30fe",
		x"10e8",
		x"60ac",
		x"00f0",
		x"10e8",
		x"00ef",
		x"10e7",
		x"00f9",
		x"40fe",
		x"10ec",
		x"00fa",
		x"a0fb",
		x"c0da",
		x"00fc",
		x"a0fb",
		x"c0da",
		x"6027",
		x"00ff",
		x"10fa",
		x"10fc",
		x"6027",
		x"0050",
		x"0048",
		x"0000",
		x"0030",
		x"0038",
		x"0004",
		x"002e",
		x"0000",
		x"0000",
		x"0017",
		x"0020",
		x"0040",
		x"0000",
		x"0040",
		x"0000",
		x"0018",
		x"0020",
		x"0018",
		x"0020",
		x"003e",
		x"003f",
		x"0001",
		x"0002",
		x"0001",
		x"0080",
		x"0003",
		x"0000",
		x"0000",
		x"0000",
		x"0003",
		x"0000",
		x"0800",
		x"0001",
		x"0000"
	);

	signal reset_counter:std_logic_vector(7 downto 0):=x"00";


	--Controls PM output to bus.
begin
	process(clk)
	begin
		if (rising_edge(clk)) then
		  bus_out <= ram(conv_integer(adress_pm));
		end if;
	end process;
	
	--Controls PM input and reset memory when button is pressed.
	process(clk)
	begin
		if (rising_edge(clk)) then
			if rst='0'then
				ram(conv_integer(reset_counter)) <= original_ram(conv_integer(reset_counter));
				reset_counter<=reset_counter+'1';
			else
				reset_counter<=x"00";
				if (pm_read = '0') then
					ram(conv_integer(adress_pm)) <= bus_in;
				end if;
			end if;
		end if;
	end process;
end Behavioral;
